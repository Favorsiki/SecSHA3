module ReOrderChiSquence(
    input [1599:0] orgin,    
    input [1599:0] reorder   
);
    assign reorder[4:0] 	= {orgin[256], orgin[192], orgin[128], orgin[64], orgin[0]};
    assign reorder[9:5] 	= {orgin[576], orgin[512], orgin[448], orgin[384], orgin[320]};
    assign reorder[14:10] 	= {orgin[896], orgin[832], orgin[768], orgin[704], orgin[640]};
    assign reorder[19:15] 	= {orgin[1216], orgin[1152], orgin[1088], orgin[1024], orgin[960]};
    assign reorder[24:20] 	= {orgin[1536], orgin[1472], orgin[1408], orgin[1344], orgin[1280]};
    assign reorder[29:25] 	= {orgin[257], orgin[193], orgin[129], orgin[65], orgin[1]};
    assign reorder[34:30] 	= {orgin[577], orgin[513], orgin[449], orgin[385], orgin[321]};
    assign reorder[39:35] 	= {orgin[897], orgin[833], orgin[769], orgin[705], orgin[641]};
    assign reorder[44:40] 	= {orgin[1217], orgin[1153], orgin[1089], orgin[1025], orgin[961]};
    assign reorder[49:45] 	= {orgin[1537], orgin[1473], orgin[1409], orgin[1345], orgin[1281]};
    assign reorder[54:50] 	= {orgin[258], orgin[194], orgin[130], orgin[66], orgin[2]};
    assign reorder[59:55] 	= {orgin[578], orgin[514], orgin[450], orgin[386], orgin[322]};
    assign reorder[64:60] 	= {orgin[898], orgin[834], orgin[770], orgin[706], orgin[642]};
    assign reorder[69:65] 	= {orgin[1218], orgin[1154], orgin[1090], orgin[1026], orgin[962]};
    assign reorder[74:70] 	= {orgin[1538], orgin[1474], orgin[1410], orgin[1346], orgin[1282]};
    assign reorder[79:75] 	= {orgin[259], orgin[195], orgin[131], orgin[67], orgin[3]};
    assign reorder[84:80] 	= {orgin[579], orgin[515], orgin[451], orgin[387], orgin[323]};
    assign reorder[89:85] 	= {orgin[899], orgin[835], orgin[771], orgin[707], orgin[643]};
    assign reorder[94:90] 	= {orgin[1219], orgin[1155], orgin[1091], orgin[1027], orgin[963]};
    assign reorder[99:95] 	= {orgin[1539], orgin[1475], orgin[1411], orgin[1347], orgin[1283]};
    assign reorder[104:100] 	= {orgin[260], orgin[196], orgin[132], orgin[68], orgin[4]};
    assign reorder[109:105] 	= {orgin[580], orgin[516], orgin[452], orgin[388], orgin[324]};
    assign reorder[114:110] 	= {orgin[900], orgin[836], orgin[772], orgin[708], orgin[644]};
    assign reorder[119:115] 	= {orgin[1220], orgin[1156], orgin[1092], orgin[1028], orgin[964]};
    assign reorder[124:120] 	= {orgin[1540], orgin[1476], orgin[1412], orgin[1348], orgin[1284]};
    assign reorder[129:125] 	= {orgin[261], orgin[197], orgin[133], orgin[69], orgin[5]};
    assign reorder[134:130] 	= {orgin[581], orgin[517], orgin[453], orgin[389], orgin[325]};
    assign reorder[139:135] 	= {orgin[901], orgin[837], orgin[773], orgin[709], orgin[645]};
    assign reorder[144:140] 	= {orgin[1221], orgin[1157], orgin[1093], orgin[1029], orgin[965]};
    assign reorder[149:145] 	= {orgin[1541], orgin[1477], orgin[1413], orgin[1349], orgin[1285]};
    assign reorder[154:150] 	= {orgin[262], orgin[198], orgin[134], orgin[70], orgin[6]};
    assign reorder[159:155] 	= {orgin[582], orgin[518], orgin[454], orgin[390], orgin[326]};
    assign reorder[164:160] 	= {orgin[902], orgin[838], orgin[774], orgin[710], orgin[646]};
    assign reorder[169:165] 	= {orgin[1222], orgin[1158], orgin[1094], orgin[1030], orgin[966]};
    assign reorder[174:170] 	= {orgin[1542], orgin[1478], orgin[1414], orgin[1350], orgin[1286]};
    assign reorder[179:175] 	= {orgin[263], orgin[199], orgin[135], orgin[71], orgin[7]};
    assign reorder[184:180] 	= {orgin[583], orgin[519], orgin[455], orgin[391], orgin[327]};
    assign reorder[189:185] 	= {orgin[903], orgin[839], orgin[775], orgin[711], orgin[647]};
    assign reorder[194:190] 	= {orgin[1223], orgin[1159], orgin[1095], orgin[1031], orgin[967]};
    assign reorder[199:195] 	= {orgin[1543], orgin[1479], orgin[1415], orgin[1351], orgin[1287]};
    assign reorder[204:200] 	= {orgin[264], orgin[200], orgin[136], orgin[72], orgin[8]};
    assign reorder[209:205] 	= {orgin[584], orgin[520], orgin[456], orgin[392], orgin[328]};
    assign reorder[214:210] 	= {orgin[904], orgin[840], orgin[776], orgin[712], orgin[648]};
    assign reorder[219:215] 	= {orgin[1224], orgin[1160], orgin[1096], orgin[1032], orgin[968]};
    assign reorder[224:220] 	= {orgin[1544], orgin[1480], orgin[1416], orgin[1352], orgin[1288]};
    assign reorder[229:225] 	= {orgin[265], orgin[201], orgin[137], orgin[73], orgin[9]};
    assign reorder[234:230] 	= {orgin[585], orgin[521], orgin[457], orgin[393], orgin[329]};
    assign reorder[239:235] 	= {orgin[905], orgin[841], orgin[777], orgin[713], orgin[649]};
    assign reorder[244:240] 	= {orgin[1225], orgin[1161], orgin[1097], orgin[1033], orgin[969]};
    assign reorder[249:245] 	= {orgin[1545], orgin[1481], orgin[1417], orgin[1353], orgin[1289]};
    assign reorder[254:250] 	= {orgin[266], orgin[202], orgin[138], orgin[74], orgin[10]};
    assign reorder[259:255] 	= {orgin[586], orgin[522], orgin[458], orgin[394], orgin[330]};
    assign reorder[264:260] 	= {orgin[906], orgin[842], orgin[778], orgin[714], orgin[650]};
    assign reorder[269:265] 	= {orgin[1226], orgin[1162], orgin[1098], orgin[1034], orgin[970]};
    assign reorder[274:270] 	= {orgin[1546], orgin[1482], orgin[1418], orgin[1354], orgin[1290]};
    assign reorder[279:275] 	= {orgin[267], orgin[203], orgin[139], orgin[75], orgin[11]};
    assign reorder[284:280] 	= {orgin[587], orgin[523], orgin[459], orgin[395], orgin[331]};
    assign reorder[289:285] 	= {orgin[907], orgin[843], orgin[779], orgin[715], orgin[651]};
    assign reorder[294:290] 	= {orgin[1227], orgin[1163], orgin[1099], orgin[1035], orgin[971]};
    assign reorder[299:295] 	= {orgin[1547], orgin[1483], orgin[1419], orgin[1355], orgin[1291]};
    assign reorder[304:300] 	= {orgin[268], orgin[204], orgin[140], orgin[76], orgin[12]};
    assign reorder[309:305] 	= {orgin[588], orgin[524], orgin[460], orgin[396], orgin[332]};
    assign reorder[314:310] 	= {orgin[908], orgin[844], orgin[780], orgin[716], orgin[652]};
    assign reorder[319:315] 	= {orgin[1228], orgin[1164], orgin[1100], orgin[1036], orgin[972]};
    assign reorder[324:320] 	= {orgin[1548], orgin[1484], orgin[1420], orgin[1356], orgin[1292]};
    assign reorder[329:325] 	= {orgin[269], orgin[205], orgin[141], orgin[77], orgin[13]};
    assign reorder[334:330] 	= {orgin[589], orgin[525], orgin[461], orgin[397], orgin[333]};
    assign reorder[339:335] 	= {orgin[909], orgin[845], orgin[781], orgin[717], orgin[653]};
    assign reorder[344:340] 	= {orgin[1229], orgin[1165], orgin[1101], orgin[1037], orgin[973]};
    assign reorder[349:345] 	= {orgin[1549], orgin[1485], orgin[1421], orgin[1357], orgin[1293]};
    assign reorder[354:350] 	= {orgin[270], orgin[206], orgin[142], orgin[78], orgin[14]};
    assign reorder[359:355] 	= {orgin[590], orgin[526], orgin[462], orgin[398], orgin[334]};
    assign reorder[364:360] 	= {orgin[910], orgin[846], orgin[782], orgin[718], orgin[654]};
    assign reorder[369:365] 	= {orgin[1230], orgin[1166], orgin[1102], orgin[1038], orgin[974]};
    assign reorder[374:370] 	= {orgin[1550], orgin[1486], orgin[1422], orgin[1358], orgin[1294]};
    assign reorder[379:375] 	= {orgin[271], orgin[207], orgin[143], orgin[79], orgin[15]};
    assign reorder[384:380] 	= {orgin[591], orgin[527], orgin[463], orgin[399], orgin[335]};
    assign reorder[389:385] 	= {orgin[911], orgin[847], orgin[783], orgin[719], orgin[655]};
    assign reorder[394:390] 	= {orgin[1231], orgin[1167], orgin[1103], orgin[1039], orgin[975]};
    assign reorder[399:395] 	= {orgin[1551], orgin[1487], orgin[1423], orgin[1359], orgin[1295]};
    assign reorder[404:400] 	= {orgin[272], orgin[208], orgin[144], orgin[80], orgin[16]};
    assign reorder[409:405] 	= {orgin[592], orgin[528], orgin[464], orgin[400], orgin[336]};
    assign reorder[414:410] 	= {orgin[912], orgin[848], orgin[784], orgin[720], orgin[656]};
    assign reorder[419:415] 	= {orgin[1232], orgin[1168], orgin[1104], orgin[1040], orgin[976]};
    assign reorder[424:420] 	= {orgin[1552], orgin[1488], orgin[1424], orgin[1360], orgin[1296]};
    assign reorder[429:425] 	= {orgin[273], orgin[209], orgin[145], orgin[81], orgin[17]};
    assign reorder[434:430] 	= {orgin[593], orgin[529], orgin[465], orgin[401], orgin[337]};
    assign reorder[439:435] 	= {orgin[913], orgin[849], orgin[785], orgin[721], orgin[657]};
    assign reorder[444:440] 	= {orgin[1233], orgin[1169], orgin[1105], orgin[1041], orgin[977]};
    assign reorder[449:445] 	= {orgin[1553], orgin[1489], orgin[1425], orgin[1361], orgin[1297]};
    assign reorder[454:450] 	= {orgin[274], orgin[210], orgin[146], orgin[82], orgin[18]};
    assign reorder[459:455] 	= {orgin[594], orgin[530], orgin[466], orgin[402], orgin[338]};
    assign reorder[464:460] 	= {orgin[914], orgin[850], orgin[786], orgin[722], orgin[658]};
    assign reorder[469:465] 	= {orgin[1234], orgin[1170], orgin[1106], orgin[1042], orgin[978]};
    assign reorder[474:470] 	= {orgin[1554], orgin[1490], orgin[1426], orgin[1362], orgin[1298]};
    assign reorder[479:475] 	= {orgin[275], orgin[211], orgin[147], orgin[83], orgin[19]};
    assign reorder[484:480] 	= {orgin[595], orgin[531], orgin[467], orgin[403], orgin[339]};
    assign reorder[489:485] 	= {orgin[915], orgin[851], orgin[787], orgin[723], orgin[659]};
    assign reorder[494:490] 	= {orgin[1235], orgin[1171], orgin[1107], orgin[1043], orgin[979]};
    assign reorder[499:495] 	= {orgin[1555], orgin[1491], orgin[1427], orgin[1363], orgin[1299]};
    assign reorder[504:500] 	= {orgin[276], orgin[212], orgin[148], orgin[84], orgin[20]};
    assign reorder[509:505] 	= {orgin[596], orgin[532], orgin[468], orgin[404], orgin[340]};
    assign reorder[514:510] 	= {orgin[916], orgin[852], orgin[788], orgin[724], orgin[660]};
    assign reorder[519:515] 	= {orgin[1236], orgin[1172], orgin[1108], orgin[1044], orgin[980]};
    assign reorder[524:520] 	= {orgin[1556], orgin[1492], orgin[1428], orgin[1364], orgin[1300]};
    assign reorder[529:525] 	= {orgin[277], orgin[213], orgin[149], orgin[85], orgin[21]};
    assign reorder[534:530] 	= {orgin[597], orgin[533], orgin[469], orgin[405], orgin[341]};
    assign reorder[539:535] 	= {orgin[917], orgin[853], orgin[789], orgin[725], orgin[661]};
    assign reorder[544:540] 	= {orgin[1237], orgin[1173], orgin[1109], orgin[1045], orgin[981]};
    assign reorder[549:545] 	= {orgin[1557], orgin[1493], orgin[1429], orgin[1365], orgin[1301]};
    assign reorder[554:550] 	= {orgin[278], orgin[214], orgin[150], orgin[86], orgin[22]};
    assign reorder[559:555] 	= {orgin[598], orgin[534], orgin[470], orgin[406], orgin[342]};
    assign reorder[564:560] 	= {orgin[918], orgin[854], orgin[790], orgin[726], orgin[662]};
    assign reorder[569:565] 	= {orgin[1238], orgin[1174], orgin[1110], orgin[1046], orgin[982]};
    assign reorder[574:570] 	= {orgin[1558], orgin[1494], orgin[1430], orgin[1366], orgin[1302]};
    assign reorder[579:575] 	= {orgin[279], orgin[215], orgin[151], orgin[87], orgin[23]};
    assign reorder[584:580] 	= {orgin[599], orgin[535], orgin[471], orgin[407], orgin[343]};
    assign reorder[589:585] 	= {orgin[919], orgin[855], orgin[791], orgin[727], orgin[663]};
    assign reorder[594:590] 	= {orgin[1239], orgin[1175], orgin[1111], orgin[1047], orgin[983]};
    assign reorder[599:595] 	= {orgin[1559], orgin[1495], orgin[1431], orgin[1367], orgin[1303]};
    assign reorder[604:600] 	= {orgin[280], orgin[216], orgin[152], orgin[88], orgin[24]};
    assign reorder[609:605] 	= {orgin[600], orgin[536], orgin[472], orgin[408], orgin[344]};
    assign reorder[614:610] 	= {orgin[920], orgin[856], orgin[792], orgin[728], orgin[664]};
    assign reorder[619:615] 	= {orgin[1240], orgin[1176], orgin[1112], orgin[1048], orgin[984]};
    assign reorder[624:620] 	= {orgin[1560], orgin[1496], orgin[1432], orgin[1368], orgin[1304]};
    assign reorder[629:625] 	= {orgin[281], orgin[217], orgin[153], orgin[89], orgin[25]};
    assign reorder[634:630] 	= {orgin[601], orgin[537], orgin[473], orgin[409], orgin[345]};
    assign reorder[639:635] 	= {orgin[921], orgin[857], orgin[793], orgin[729], orgin[665]};
    assign reorder[644:640] 	= {orgin[1241], orgin[1177], orgin[1113], orgin[1049], orgin[985]};
    assign reorder[649:645] 	= {orgin[1561], orgin[1497], orgin[1433], orgin[1369], orgin[1305]};
    assign reorder[654:650] 	= {orgin[282], orgin[218], orgin[154], orgin[90], orgin[26]};
    assign reorder[659:655] 	= {orgin[602], orgin[538], orgin[474], orgin[410], orgin[346]};
    assign reorder[664:660] 	= {orgin[922], orgin[858], orgin[794], orgin[730], orgin[666]};
    assign reorder[669:665] 	= {orgin[1242], orgin[1178], orgin[1114], orgin[1050], orgin[986]};
    assign reorder[674:670] 	= {orgin[1562], orgin[1498], orgin[1434], orgin[1370], orgin[1306]};
    assign reorder[679:675] 	= {orgin[283], orgin[219], orgin[155], orgin[91], orgin[27]};
    assign reorder[684:680] 	= {orgin[603], orgin[539], orgin[475], orgin[411], orgin[347]};
    assign reorder[689:685] 	= {orgin[923], orgin[859], orgin[795], orgin[731], orgin[667]};
    assign reorder[694:690] 	= {orgin[1243], orgin[1179], orgin[1115], orgin[1051], orgin[987]};
    assign reorder[699:695] 	= {orgin[1563], orgin[1499], orgin[1435], orgin[1371], orgin[1307]};
    assign reorder[704:700] 	= {orgin[284], orgin[220], orgin[156], orgin[92], orgin[28]};
    assign reorder[709:705] 	= {orgin[604], orgin[540], orgin[476], orgin[412], orgin[348]};
    assign reorder[714:710] 	= {orgin[924], orgin[860], orgin[796], orgin[732], orgin[668]};
    assign reorder[719:715] 	= {orgin[1244], orgin[1180], orgin[1116], orgin[1052], orgin[988]};
    assign reorder[724:720] 	= {orgin[1564], orgin[1500], orgin[1436], orgin[1372], orgin[1308]};
    assign reorder[729:725] 	= {orgin[285], orgin[221], orgin[157], orgin[93], orgin[29]};
    assign reorder[734:730] 	= {orgin[605], orgin[541], orgin[477], orgin[413], orgin[349]};
    assign reorder[739:735] 	= {orgin[925], orgin[861], orgin[797], orgin[733], orgin[669]};
    assign reorder[744:740] 	= {orgin[1245], orgin[1181], orgin[1117], orgin[1053], orgin[989]};
    assign reorder[749:745] 	= {orgin[1565], orgin[1501], orgin[1437], orgin[1373], orgin[1309]};
    assign reorder[754:750] 	= {orgin[286], orgin[222], orgin[158], orgin[94], orgin[30]};
    assign reorder[759:755] 	= {orgin[606], orgin[542], orgin[478], orgin[414], orgin[350]};
    assign reorder[764:760] 	= {orgin[926], orgin[862], orgin[798], orgin[734], orgin[670]};
    assign reorder[769:765] 	= {orgin[1246], orgin[1182], orgin[1118], orgin[1054], orgin[990]};
    assign reorder[774:770] 	= {orgin[1566], orgin[1502], orgin[1438], orgin[1374], orgin[1310]};
    assign reorder[779:775] 	= {orgin[287], orgin[223], orgin[159], orgin[95], orgin[31]};
    assign reorder[784:780] 	= {orgin[607], orgin[543], orgin[479], orgin[415], orgin[351]};
    assign reorder[789:785] 	= {orgin[927], orgin[863], orgin[799], orgin[735], orgin[671]};
    assign reorder[794:790] 	= {orgin[1247], orgin[1183], orgin[1119], orgin[1055], orgin[991]};
    assign reorder[799:795] 	= {orgin[1567], orgin[1503], orgin[1439], orgin[1375], orgin[1311]};
    assign reorder[804:800] 	= {orgin[288], orgin[224], orgin[160], orgin[96], orgin[32]};
    assign reorder[809:805] 	= {orgin[608], orgin[544], orgin[480], orgin[416], orgin[352]};
    assign reorder[814:810] 	= {orgin[928], orgin[864], orgin[800], orgin[736], orgin[672]};
    assign reorder[819:815] 	= {orgin[1248], orgin[1184], orgin[1120], orgin[1056], orgin[992]};
    assign reorder[824:820] 	= {orgin[1568], orgin[1504], orgin[1440], orgin[1376], orgin[1312]};
    assign reorder[829:825] 	= {orgin[289], orgin[225], orgin[161], orgin[97], orgin[33]};
    assign reorder[834:830] 	= {orgin[609], orgin[545], orgin[481], orgin[417], orgin[353]};
    assign reorder[839:835] 	= {orgin[929], orgin[865], orgin[801], orgin[737], orgin[673]};
    assign reorder[844:840] 	= {orgin[1249], orgin[1185], orgin[1121], orgin[1057], orgin[993]};
    assign reorder[849:845] 	= {orgin[1569], orgin[1505], orgin[1441], orgin[1377], orgin[1313]};
    assign reorder[854:850] 	= {orgin[290], orgin[226], orgin[162], orgin[98], orgin[34]};
    assign reorder[859:855] 	= {orgin[610], orgin[546], orgin[482], orgin[418], orgin[354]};
    assign reorder[864:860] 	= {orgin[930], orgin[866], orgin[802], orgin[738], orgin[674]};
    assign reorder[869:865] 	= {orgin[1250], orgin[1186], orgin[1122], orgin[1058], orgin[994]};
    assign reorder[874:870] 	= {orgin[1570], orgin[1506], orgin[1442], orgin[1378], orgin[1314]};
    assign reorder[879:875] 	= {orgin[291], orgin[227], orgin[163], orgin[99], orgin[35]};
    assign reorder[884:880] 	= {orgin[611], orgin[547], orgin[483], orgin[419], orgin[355]};
    assign reorder[889:885] 	= {orgin[931], orgin[867], orgin[803], orgin[739], orgin[675]};
    assign reorder[894:890] 	= {orgin[1251], orgin[1187], orgin[1123], orgin[1059], orgin[995]};
    assign reorder[899:895] 	= {orgin[1571], orgin[1507], orgin[1443], orgin[1379], orgin[1315]};
    assign reorder[904:900] 	= {orgin[292], orgin[228], orgin[164], orgin[100], orgin[36]};
    assign reorder[909:905] 	= {orgin[612], orgin[548], orgin[484], orgin[420], orgin[356]};
    assign reorder[914:910] 	= {orgin[932], orgin[868], orgin[804], orgin[740], orgin[676]};
    assign reorder[919:915] 	= {orgin[1252], orgin[1188], orgin[1124], orgin[1060], orgin[996]};
    assign reorder[924:920] 	= {orgin[1572], orgin[1508], orgin[1444], orgin[1380], orgin[1316]};
    assign reorder[929:925] 	= {orgin[293], orgin[229], orgin[165], orgin[101], orgin[37]};
    assign reorder[934:930] 	= {orgin[613], orgin[549], orgin[485], orgin[421], orgin[357]};
    assign reorder[939:935] 	= {orgin[933], orgin[869], orgin[805], orgin[741], orgin[677]};
    assign reorder[944:940] 	= {orgin[1253], orgin[1189], orgin[1125], orgin[1061], orgin[997]};
    assign reorder[949:945] 	= {orgin[1573], orgin[1509], orgin[1445], orgin[1381], orgin[1317]};
    assign reorder[954:950] 	= {orgin[294], orgin[230], orgin[166], orgin[102], orgin[38]};
    assign reorder[959:955] 	= {orgin[614], orgin[550], orgin[486], orgin[422], orgin[358]};
    assign reorder[964:960] 	= {orgin[934], orgin[870], orgin[806], orgin[742], orgin[678]};
    assign reorder[969:965] 	= {orgin[1254], orgin[1190], orgin[1126], orgin[1062], orgin[998]};
    assign reorder[974:970] 	= {orgin[1574], orgin[1510], orgin[1446], orgin[1382], orgin[1318]};
    assign reorder[979:975] 	= {orgin[295], orgin[231], orgin[167], orgin[103], orgin[39]};
    assign reorder[984:980] 	= {orgin[615], orgin[551], orgin[487], orgin[423], orgin[359]};
    assign reorder[989:985] 	= {orgin[935], orgin[871], orgin[807], orgin[743], orgin[679]};
    assign reorder[994:990] 	= {orgin[1255], orgin[1191], orgin[1127], orgin[1063], orgin[999]};
    assign reorder[999:995] 	= {orgin[1575], orgin[1511], orgin[1447], orgin[1383], orgin[1319]};
    assign reorder[1004:1000] 	= {orgin[296], orgin[232], orgin[168], orgin[104], orgin[40]};
    assign reorder[1009:1005] 	= {orgin[616], orgin[552], orgin[488], orgin[424], orgin[360]};
    assign reorder[1014:1010] 	= {orgin[936], orgin[872], orgin[808], orgin[744], orgin[680]};
    assign reorder[1019:1015] 	= {orgin[1256], orgin[1192], orgin[1128], orgin[1064], orgin[1000]};
    assign reorder[1024:1020] 	= {orgin[1576], orgin[1512], orgin[1448], orgin[1384], orgin[1320]};
    assign reorder[1029:1025] 	= {orgin[297], orgin[233], orgin[169], orgin[105], orgin[41]};
    assign reorder[1034:1030] 	= {orgin[617], orgin[553], orgin[489], orgin[425], orgin[361]};
    assign reorder[1039:1035] 	= {orgin[937], orgin[873], orgin[809], orgin[745], orgin[681]};
    assign reorder[1044:1040] 	= {orgin[1257], orgin[1193], orgin[1129], orgin[1065], orgin[1001]};
    assign reorder[1049:1045] 	= {orgin[1577], orgin[1513], orgin[1449], orgin[1385], orgin[1321]};
    assign reorder[1054:1050] 	= {orgin[298], orgin[234], orgin[170], orgin[106], orgin[42]};
    assign reorder[1059:1055] 	= {orgin[618], orgin[554], orgin[490], orgin[426], orgin[362]};
    assign reorder[1064:1060] 	= {orgin[938], orgin[874], orgin[810], orgin[746], orgin[682]};
    assign reorder[1069:1065] 	= {orgin[1258], orgin[1194], orgin[1130], orgin[1066], orgin[1002]};
    assign reorder[1074:1070] 	= {orgin[1578], orgin[1514], orgin[1450], orgin[1386], orgin[1322]};
    assign reorder[1079:1075] 	= {orgin[299], orgin[235], orgin[171], orgin[107], orgin[43]};
    assign reorder[1084:1080] 	= {orgin[619], orgin[555], orgin[491], orgin[427], orgin[363]};
    assign reorder[1089:1085] 	= {orgin[939], orgin[875], orgin[811], orgin[747], orgin[683]};
    assign reorder[1094:1090] 	= {orgin[1259], orgin[1195], orgin[1131], orgin[1067], orgin[1003]};
    assign reorder[1099:1095] 	= {orgin[1579], orgin[1515], orgin[1451], orgin[1387], orgin[1323]};
    assign reorder[1104:1100] 	= {orgin[300], orgin[236], orgin[172], orgin[108], orgin[44]};
    assign reorder[1109:1105] 	= {orgin[620], orgin[556], orgin[492], orgin[428], orgin[364]};
    assign reorder[1114:1110] 	= {orgin[940], orgin[876], orgin[812], orgin[748], orgin[684]};
    assign reorder[1119:1115] 	= {orgin[1260], orgin[1196], orgin[1132], orgin[1068], orgin[1004]};
    assign reorder[1124:1120] 	= {orgin[1580], orgin[1516], orgin[1452], orgin[1388], orgin[1324]};
    assign reorder[1129:1125] 	= {orgin[301], orgin[237], orgin[173], orgin[109], orgin[45]};
    assign reorder[1134:1130] 	= {orgin[621], orgin[557], orgin[493], orgin[429], orgin[365]};
    assign reorder[1139:1135] 	= {orgin[941], orgin[877], orgin[813], orgin[749], orgin[685]};
    assign reorder[1144:1140] 	= {orgin[1261], orgin[1197], orgin[1133], orgin[1069], orgin[1005]};
    assign reorder[1149:1145] 	= {orgin[1581], orgin[1517], orgin[1453], orgin[1389], orgin[1325]};
    assign reorder[1154:1150] 	= {orgin[302], orgin[238], orgin[174], orgin[110], orgin[46]};
    assign reorder[1159:1155] 	= {orgin[622], orgin[558], orgin[494], orgin[430], orgin[366]};
    assign reorder[1164:1160] 	= {orgin[942], orgin[878], orgin[814], orgin[750], orgin[686]};
    assign reorder[1169:1165] 	= {orgin[1262], orgin[1198], orgin[1134], orgin[1070], orgin[1006]};
    assign reorder[1174:1170] 	= {orgin[1582], orgin[1518], orgin[1454], orgin[1390], orgin[1326]};
    assign reorder[1179:1175] 	= {orgin[303], orgin[239], orgin[175], orgin[111], orgin[47]};
    assign reorder[1184:1180] 	= {orgin[623], orgin[559], orgin[495], orgin[431], orgin[367]};
    assign reorder[1189:1185] 	= {orgin[943], orgin[879], orgin[815], orgin[751], orgin[687]};
    assign reorder[1194:1190] 	= {orgin[1263], orgin[1199], orgin[1135], orgin[1071], orgin[1007]};
    assign reorder[1199:1195] 	= {orgin[1583], orgin[1519], orgin[1455], orgin[1391], orgin[1327]};
    assign reorder[1204:1200] 	= {orgin[304], orgin[240], orgin[176], orgin[112], orgin[48]};
    assign reorder[1209:1205] 	= {orgin[624], orgin[560], orgin[496], orgin[432], orgin[368]};
    assign reorder[1214:1210] 	= {orgin[944], orgin[880], orgin[816], orgin[752], orgin[688]};
    assign reorder[1219:1215] 	= {orgin[1264], orgin[1200], orgin[1136], orgin[1072], orgin[1008]};
    assign reorder[1224:1220] 	= {orgin[1584], orgin[1520], orgin[1456], orgin[1392], orgin[1328]};
    assign reorder[1229:1225] 	= {orgin[305], orgin[241], orgin[177], orgin[113], orgin[49]};
    assign reorder[1234:1230] 	= {orgin[625], orgin[561], orgin[497], orgin[433], orgin[369]};
    assign reorder[1239:1235] 	= {orgin[945], orgin[881], orgin[817], orgin[753], orgin[689]};
    assign reorder[1244:1240] 	= {orgin[1265], orgin[1201], orgin[1137], orgin[1073], orgin[1009]};
    assign reorder[1249:1245] 	= {orgin[1585], orgin[1521], orgin[1457], orgin[1393], orgin[1329]};
    assign reorder[1254:1250] 	= {orgin[306], orgin[242], orgin[178], orgin[114], orgin[50]};
    assign reorder[1259:1255] 	= {orgin[626], orgin[562], orgin[498], orgin[434], orgin[370]};
    assign reorder[1264:1260] 	= {orgin[946], orgin[882], orgin[818], orgin[754], orgin[690]};
    assign reorder[1269:1265] 	= {orgin[1266], orgin[1202], orgin[1138], orgin[1074], orgin[1010]};
    assign reorder[1274:1270] 	= {orgin[1586], orgin[1522], orgin[1458], orgin[1394], orgin[1330]};
    assign reorder[1279:1275] 	= {orgin[307], orgin[243], orgin[179], orgin[115], orgin[51]};
    assign reorder[1284:1280] 	= {orgin[627], orgin[563], orgin[499], orgin[435], orgin[371]};
    assign reorder[1289:1285] 	= {orgin[947], orgin[883], orgin[819], orgin[755], orgin[691]};
    assign reorder[1294:1290] 	= {orgin[1267], orgin[1203], orgin[1139], orgin[1075], orgin[1011]};
    assign reorder[1299:1295] 	= {orgin[1587], orgin[1523], orgin[1459], orgin[1395], orgin[1331]};
    assign reorder[1304:1300] 	= {orgin[308], orgin[244], orgin[180], orgin[116], orgin[52]};
    assign reorder[1309:1305] 	= {orgin[628], orgin[564], orgin[500], orgin[436], orgin[372]};
    assign reorder[1314:1310] 	= {orgin[948], orgin[884], orgin[820], orgin[756], orgin[692]};
    assign reorder[1319:1315] 	= {orgin[1268], orgin[1204], orgin[1140], orgin[1076], orgin[1012]};
    assign reorder[1324:1320] 	= {orgin[1588], orgin[1524], orgin[1460], orgin[1396], orgin[1332]};
    assign reorder[1329:1325] 	= {orgin[309], orgin[245], orgin[181], orgin[117], orgin[53]};
    assign reorder[1334:1330] 	= {orgin[629], orgin[565], orgin[501], orgin[437], orgin[373]};
    assign reorder[1339:1335] 	= {orgin[949], orgin[885], orgin[821], orgin[757], orgin[693]};
    assign reorder[1344:1340] 	= {orgin[1269], orgin[1205], orgin[1141], orgin[1077], orgin[1013]};
    assign reorder[1349:1345] 	= {orgin[1589], orgin[1525], orgin[1461], orgin[1397], orgin[1333]};
    assign reorder[1354:1350] 	= {orgin[310], orgin[246], orgin[182], orgin[118], orgin[54]};
    assign reorder[1359:1355] 	= {orgin[630], orgin[566], orgin[502], orgin[438], orgin[374]};
    assign reorder[1364:1360] 	= {orgin[950], orgin[886], orgin[822], orgin[758], orgin[694]};
    assign reorder[1369:1365] 	= {orgin[1270], orgin[1206], orgin[1142], orgin[1078], orgin[1014]};
    assign reorder[1374:1370] 	= {orgin[1590], orgin[1526], orgin[1462], orgin[1398], orgin[1334]};
    assign reorder[1379:1375] 	= {orgin[311], orgin[247], orgin[183], orgin[119], orgin[55]};
    assign reorder[1384:1380] 	= {orgin[631], orgin[567], orgin[503], orgin[439], orgin[375]};
    assign reorder[1389:1385] 	= {orgin[951], orgin[887], orgin[823], orgin[759], orgin[695]};
    assign reorder[1394:1390] 	= {orgin[1271], orgin[1207], orgin[1143], orgin[1079], orgin[1015]};
    assign reorder[1399:1395] 	= {orgin[1591], orgin[1527], orgin[1463], orgin[1399], orgin[1335]};
    assign reorder[1404:1400] 	= {orgin[312], orgin[248], orgin[184], orgin[120], orgin[56]};
    assign reorder[1409:1405] 	= {orgin[632], orgin[568], orgin[504], orgin[440], orgin[376]};
    assign reorder[1414:1410] 	= {orgin[952], orgin[888], orgin[824], orgin[760], orgin[696]};
    assign reorder[1419:1415] 	= {orgin[1272], orgin[1208], orgin[1144], orgin[1080], orgin[1016]};
    assign reorder[1424:1420] 	= {orgin[1592], orgin[1528], orgin[1464], orgin[1400], orgin[1336]};
    assign reorder[1429:1425] 	= {orgin[313], orgin[249], orgin[185], orgin[121], orgin[57]};
    assign reorder[1434:1430] 	= {orgin[633], orgin[569], orgin[505], orgin[441], orgin[377]};
    assign reorder[1439:1435] 	= {orgin[953], orgin[889], orgin[825], orgin[761], orgin[697]};
    assign reorder[1444:1440] 	= {orgin[1273], orgin[1209], orgin[1145], orgin[1081], orgin[1017]};
    assign reorder[1449:1445] 	= {orgin[1593], orgin[1529], orgin[1465], orgin[1401], orgin[1337]};
    assign reorder[1454:1450] 	= {orgin[314], orgin[250], orgin[186], orgin[122], orgin[58]};
    assign reorder[1459:1455] 	= {orgin[634], orgin[570], orgin[506], orgin[442], orgin[378]};
    assign reorder[1464:1460] 	= {orgin[954], orgin[890], orgin[826], orgin[762], orgin[698]};
    assign reorder[1469:1465] 	= {orgin[1274], orgin[1210], orgin[1146], orgin[1082], orgin[1018]};
    assign reorder[1474:1470] 	= {orgin[1594], orgin[1530], orgin[1466], orgin[1402], orgin[1338]};
    assign reorder[1479:1475] 	= {orgin[315], orgin[251], orgin[187], orgin[123], orgin[59]};
    assign reorder[1484:1480] 	= {orgin[635], orgin[571], orgin[507], orgin[443], orgin[379]};
    assign reorder[1489:1485] 	= {orgin[955], orgin[891], orgin[827], orgin[763], orgin[699]};
    assign reorder[1494:1490] 	= {orgin[1275], orgin[1211], orgin[1147], orgin[1083], orgin[1019]};
    assign reorder[1499:1495] 	= {orgin[1595], orgin[1531], orgin[1467], orgin[1403], orgin[1339]};
    assign reorder[1504:1500] 	= {orgin[316], orgin[252], orgin[188], orgin[124], orgin[60]};
    assign reorder[1509:1505] 	= {orgin[636], orgin[572], orgin[508], orgin[444], orgin[380]};
    assign reorder[1514:1510] 	= {orgin[956], orgin[892], orgin[828], orgin[764], orgin[700]};
    assign reorder[1519:1515] 	= {orgin[1276], orgin[1212], orgin[1148], orgin[1084], orgin[1020]};
    assign reorder[1524:1520] 	= {orgin[1596], orgin[1532], orgin[1468], orgin[1404], orgin[1340]};
    assign reorder[1529:1525] 	= {orgin[317], orgin[253], orgin[189], orgin[125], orgin[61]};
    assign reorder[1534:1530] 	= {orgin[637], orgin[573], orgin[509], orgin[445], orgin[381]};
    assign reorder[1539:1535] 	= {orgin[957], orgin[893], orgin[829], orgin[765], orgin[701]};
    assign reorder[1544:1540] 	= {orgin[1277], orgin[1213], orgin[1149], orgin[1085], orgin[1021]};
    assign reorder[1549:1545] 	= {orgin[1597], orgin[1533], orgin[1469], orgin[1405], orgin[1341]};
    assign reorder[1554:1550] 	= {orgin[318], orgin[254], orgin[190], orgin[126], orgin[62]};
    assign reorder[1559:1555] 	= {orgin[638], orgin[574], orgin[510], orgin[446], orgin[382]};
    assign reorder[1564:1560] 	= {orgin[958], orgin[894], orgin[830], orgin[766], orgin[702]};
    assign reorder[1569:1565] 	= {orgin[1278], orgin[1214], orgin[1150], orgin[1086], orgin[1022]};
    assign reorder[1574:1570] 	= {orgin[1598], orgin[1534], orgin[1470], orgin[1406], orgin[1342]};
    assign reorder[1579:1575] 	= {orgin[319], orgin[255], orgin[191], orgin[127], orgin[63]};
    assign reorder[1584:1580] 	= {orgin[639], orgin[575], orgin[511], orgin[447], orgin[383]};
    assign reorder[1589:1585] 	= {orgin[959], orgin[895], orgin[831], orgin[767], orgin[703]};
    assign reorder[1594:1590] 	= {orgin[1279], orgin[1215], orgin[1151], orgin[1087], orgin[1023]};
    assign reorder[1599:1595] 	= {orgin[1599], orgin[1535], orgin[1471], orgin[1407], orgin[1343]};
endmodule


module InvReOrderChiSquence(
    input [1599:0] reorder,    
    input [1599:0] orgin     
);
    assign {orgin[256], orgin[192], orgin[128], orgin[64], orgin[0]} 	= reorder[4:0];
    assign {orgin[576], orgin[512], orgin[448], orgin[384], orgin[320]} 	= reorder[9:5];
    assign {orgin[896], orgin[832], orgin[768], orgin[704], orgin[640]} 	= reorder[14:10];
    assign {orgin[1216], orgin[1152], orgin[1088], orgin[1024], orgin[960]} 	= reorder[19:15];
    assign {orgin[1536], orgin[1472], orgin[1408], orgin[1344], orgin[1280]} 	= reorder[24:20];
    assign {orgin[257], orgin[193], orgin[129], orgin[65], orgin[1]} 	= reorder[29:25];
    assign {orgin[577], orgin[513], orgin[449], orgin[385], orgin[321]} 	= reorder[34:30];
    assign {orgin[897], orgin[833], orgin[769], orgin[705], orgin[641]} 	= reorder[39:35];
    assign {orgin[1217], orgin[1153], orgin[1089], orgin[1025], orgin[961]} 	= reorder[44:40];
    assign {orgin[1537], orgin[1473], orgin[1409], orgin[1345], orgin[1281]} 	= reorder[49:45];
    assign {orgin[258], orgin[194], orgin[130], orgin[66], orgin[2]} 	= reorder[54:50];
    assign {orgin[578], orgin[514], orgin[450], orgin[386], orgin[322]} 	= reorder[59:55];
    assign {orgin[898], orgin[834], orgin[770], orgin[706], orgin[642]} 	= reorder[64:60];
    assign {orgin[1218], orgin[1154], orgin[1090], orgin[1026], orgin[962]} 	= reorder[69:65];
    assign {orgin[1538], orgin[1474], orgin[1410], orgin[1346], orgin[1282]} 	= reorder[74:70];
    assign {orgin[259], orgin[195], orgin[131], orgin[67], orgin[3]} 	= reorder[79:75];
    assign {orgin[579], orgin[515], orgin[451], orgin[387], orgin[323]} 	= reorder[84:80];
    assign {orgin[899], orgin[835], orgin[771], orgin[707], orgin[643]} 	= reorder[89:85];
    assign {orgin[1219], orgin[1155], orgin[1091], orgin[1027], orgin[963]} 	= reorder[94:90];
    assign {orgin[1539], orgin[1475], orgin[1411], orgin[1347], orgin[1283]} 	= reorder[99:95];
    assign {orgin[260], orgin[196], orgin[132], orgin[68], orgin[4]} 	= reorder[104:100];
    assign {orgin[580], orgin[516], orgin[452], orgin[388], orgin[324]} 	= reorder[109:105];
    assign {orgin[900], orgin[836], orgin[772], orgin[708], orgin[644]} 	= reorder[114:110];
    assign {orgin[1220], orgin[1156], orgin[1092], orgin[1028], orgin[964]} 	= reorder[119:115];
    assign {orgin[1540], orgin[1476], orgin[1412], orgin[1348], orgin[1284]} 	= reorder[124:120];
    assign {orgin[261], orgin[197], orgin[133], orgin[69], orgin[5]} 	= reorder[129:125];
    assign {orgin[581], orgin[517], orgin[453], orgin[389], orgin[325]} 	= reorder[134:130];
    assign {orgin[901], orgin[837], orgin[773], orgin[709], orgin[645]} 	= reorder[139:135];
    assign {orgin[1221], orgin[1157], orgin[1093], orgin[1029], orgin[965]} 	= reorder[144:140];
    assign {orgin[1541], orgin[1477], orgin[1413], orgin[1349], orgin[1285]} 	= reorder[149:145];
    assign {orgin[262], orgin[198], orgin[134], orgin[70], orgin[6]} 	= reorder[154:150];
    assign {orgin[582], orgin[518], orgin[454], orgin[390], orgin[326]} 	= reorder[159:155];
    assign {orgin[902], orgin[838], orgin[774], orgin[710], orgin[646]} 	= reorder[164:160];
    assign {orgin[1222], orgin[1158], orgin[1094], orgin[1030], orgin[966]} 	= reorder[169:165];
    assign {orgin[1542], orgin[1478], orgin[1414], orgin[1350], orgin[1286]} 	= reorder[174:170];
    assign {orgin[263], orgin[199], orgin[135], orgin[71], orgin[7]} 	= reorder[179:175];
    assign {orgin[583], orgin[519], orgin[455], orgin[391], orgin[327]} 	= reorder[184:180];
    assign {orgin[903], orgin[839], orgin[775], orgin[711], orgin[647]} 	= reorder[189:185];
    assign {orgin[1223], orgin[1159], orgin[1095], orgin[1031], orgin[967]} 	= reorder[194:190];
    assign {orgin[1543], orgin[1479], orgin[1415], orgin[1351], orgin[1287]} 	= reorder[199:195];
    assign {orgin[264], orgin[200], orgin[136], orgin[72], orgin[8]} 	= reorder[204:200];
    assign {orgin[584], orgin[520], orgin[456], orgin[392], orgin[328]} 	= reorder[209:205];
    assign {orgin[904], orgin[840], orgin[776], orgin[712], orgin[648]} 	= reorder[214:210];
    assign {orgin[1224], orgin[1160], orgin[1096], orgin[1032], orgin[968]} 	= reorder[219:215];
    assign {orgin[1544], orgin[1480], orgin[1416], orgin[1352], orgin[1288]} 	= reorder[224:220];
    assign {orgin[265], orgin[201], orgin[137], orgin[73], orgin[9]} 	= reorder[229:225];
    assign {orgin[585], orgin[521], orgin[457], orgin[393], orgin[329]} 	= reorder[234:230];
    assign {orgin[905], orgin[841], orgin[777], orgin[713], orgin[649]} 	= reorder[239:235];
    assign {orgin[1225], orgin[1161], orgin[1097], orgin[1033], orgin[969]} 	= reorder[244:240];
    assign {orgin[1545], orgin[1481], orgin[1417], orgin[1353], orgin[1289]} 	= reorder[249:245];
    assign {orgin[266], orgin[202], orgin[138], orgin[74], orgin[10]} 	= reorder[254:250];
    assign {orgin[586], orgin[522], orgin[458], orgin[394], orgin[330]} 	= reorder[259:255];
    assign {orgin[906], orgin[842], orgin[778], orgin[714], orgin[650]} 	= reorder[264:260];
    assign {orgin[1226], orgin[1162], orgin[1098], orgin[1034], orgin[970]} 	= reorder[269:265];
    assign {orgin[1546], orgin[1482], orgin[1418], orgin[1354], orgin[1290]} 	= reorder[274:270];
    assign {orgin[267], orgin[203], orgin[139], orgin[75], orgin[11]} 	= reorder[279:275];
    assign {orgin[587], orgin[523], orgin[459], orgin[395], orgin[331]} 	= reorder[284:280];
    assign {orgin[907], orgin[843], orgin[779], orgin[715], orgin[651]} 	= reorder[289:285];
    assign {orgin[1227], orgin[1163], orgin[1099], orgin[1035], orgin[971]} 	= reorder[294:290];
    assign {orgin[1547], orgin[1483], orgin[1419], orgin[1355], orgin[1291]} 	= reorder[299:295];
    assign {orgin[268], orgin[204], orgin[140], orgin[76], orgin[12]} 	= reorder[304:300];
    assign {orgin[588], orgin[524], orgin[460], orgin[396], orgin[332]} 	= reorder[309:305];
    assign {orgin[908], orgin[844], orgin[780], orgin[716], orgin[652]} 	= reorder[314:310];
    assign {orgin[1228], orgin[1164], orgin[1100], orgin[1036], orgin[972]} 	= reorder[319:315];
    assign {orgin[1548], orgin[1484], orgin[1420], orgin[1356], orgin[1292]} 	= reorder[324:320];
    assign {orgin[269], orgin[205], orgin[141], orgin[77], orgin[13]} 	= reorder[329:325];
    assign {orgin[589], orgin[525], orgin[461], orgin[397], orgin[333]} 	= reorder[334:330];
    assign {orgin[909], orgin[845], orgin[781], orgin[717], orgin[653]} 	= reorder[339:335];
    assign {orgin[1229], orgin[1165], orgin[1101], orgin[1037], orgin[973]} 	= reorder[344:340];
    assign {orgin[1549], orgin[1485], orgin[1421], orgin[1357], orgin[1293]} 	= reorder[349:345];
    assign {orgin[270], orgin[206], orgin[142], orgin[78], orgin[14]} 	= reorder[354:350];
    assign {orgin[590], orgin[526], orgin[462], orgin[398], orgin[334]} 	= reorder[359:355];
    assign {orgin[910], orgin[846], orgin[782], orgin[718], orgin[654]} 	= reorder[364:360];
    assign {orgin[1230], orgin[1166], orgin[1102], orgin[1038], orgin[974]} 	= reorder[369:365];
    assign {orgin[1550], orgin[1486], orgin[1422], orgin[1358], orgin[1294]} 	= reorder[374:370];
    assign {orgin[271], orgin[207], orgin[143], orgin[79], orgin[15]} 	= reorder[379:375];
    assign {orgin[591], orgin[527], orgin[463], orgin[399], orgin[335]} 	= reorder[384:380];
    assign {orgin[911], orgin[847], orgin[783], orgin[719], orgin[655]} 	= reorder[389:385];
    assign {orgin[1231], orgin[1167], orgin[1103], orgin[1039], orgin[975]} 	= reorder[394:390];
    assign {orgin[1551], orgin[1487], orgin[1423], orgin[1359], orgin[1295]} 	= reorder[399:395];
    assign {orgin[272], orgin[208], orgin[144], orgin[80], orgin[16]} 	= reorder[404:400];
    assign {orgin[592], orgin[528], orgin[464], orgin[400], orgin[336]} 	= reorder[409:405];
    assign {orgin[912], orgin[848], orgin[784], orgin[720], orgin[656]} 	= reorder[414:410];
    assign {orgin[1232], orgin[1168], orgin[1104], orgin[1040], orgin[976]} 	= reorder[419:415];
    assign {orgin[1552], orgin[1488], orgin[1424], orgin[1360], orgin[1296]} 	= reorder[424:420];
    assign {orgin[273], orgin[209], orgin[145], orgin[81], orgin[17]} 	= reorder[429:425];
    assign {orgin[593], orgin[529], orgin[465], orgin[401], orgin[337]} 	= reorder[434:430];
    assign {orgin[913], orgin[849], orgin[785], orgin[721], orgin[657]} 	= reorder[439:435];
    assign {orgin[1233], orgin[1169], orgin[1105], orgin[1041], orgin[977]} 	= reorder[444:440];
    assign {orgin[1553], orgin[1489], orgin[1425], orgin[1361], orgin[1297]} 	= reorder[449:445];
    assign {orgin[274], orgin[210], orgin[146], orgin[82], orgin[18]} 	= reorder[454:450];
    assign {orgin[594], orgin[530], orgin[466], orgin[402], orgin[338]} 	= reorder[459:455];
    assign {orgin[914], orgin[850], orgin[786], orgin[722], orgin[658]} 	= reorder[464:460];
    assign {orgin[1234], orgin[1170], orgin[1106], orgin[1042], orgin[978]} 	= reorder[469:465];
    assign {orgin[1554], orgin[1490], orgin[1426], orgin[1362], orgin[1298]} 	= reorder[474:470];
    assign {orgin[275], orgin[211], orgin[147], orgin[83], orgin[19]} 	= reorder[479:475];
    assign {orgin[595], orgin[531], orgin[467], orgin[403], orgin[339]} 	= reorder[484:480];
    assign {orgin[915], orgin[851], orgin[787], orgin[723], orgin[659]} 	= reorder[489:485];
    assign {orgin[1235], orgin[1171], orgin[1107], orgin[1043], orgin[979]} 	= reorder[494:490];
    assign {orgin[1555], orgin[1491], orgin[1427], orgin[1363], orgin[1299]} 	= reorder[499:495];
    assign {orgin[276], orgin[212], orgin[148], orgin[84], orgin[20]} 	= reorder[504:500];
    assign {orgin[596], orgin[532], orgin[468], orgin[404], orgin[340]} 	= reorder[509:505];
    assign {orgin[916], orgin[852], orgin[788], orgin[724], orgin[660]} 	= reorder[514:510];
    assign {orgin[1236], orgin[1172], orgin[1108], orgin[1044], orgin[980]} 	= reorder[519:515];
    assign {orgin[1556], orgin[1492], orgin[1428], orgin[1364], orgin[1300]} 	= reorder[524:520];
    assign {orgin[277], orgin[213], orgin[149], orgin[85], orgin[21]} 	= reorder[529:525];
    assign {orgin[597], orgin[533], orgin[469], orgin[405], orgin[341]} 	= reorder[534:530];
    assign {orgin[917], orgin[853], orgin[789], orgin[725], orgin[661]} 	= reorder[539:535];
    assign {orgin[1237], orgin[1173], orgin[1109], orgin[1045], orgin[981]} 	= reorder[544:540];
    assign {orgin[1557], orgin[1493], orgin[1429], orgin[1365], orgin[1301]} 	= reorder[549:545];
    assign {orgin[278], orgin[214], orgin[150], orgin[86], orgin[22]} 	= reorder[554:550];
    assign {orgin[598], orgin[534], orgin[470], orgin[406], orgin[342]} 	= reorder[559:555];
    assign {orgin[918], orgin[854], orgin[790], orgin[726], orgin[662]} 	= reorder[564:560];
    assign {orgin[1238], orgin[1174], orgin[1110], orgin[1046], orgin[982]} 	= reorder[569:565];
    assign {orgin[1558], orgin[1494], orgin[1430], orgin[1366], orgin[1302]} 	= reorder[574:570];
    assign {orgin[279], orgin[215], orgin[151], orgin[87], orgin[23]} 	= reorder[579:575];
    assign {orgin[599], orgin[535], orgin[471], orgin[407], orgin[343]} 	= reorder[584:580];
    assign {orgin[919], orgin[855], orgin[791], orgin[727], orgin[663]} 	= reorder[589:585];
    assign {orgin[1239], orgin[1175], orgin[1111], orgin[1047], orgin[983]} 	= reorder[594:590];
    assign {orgin[1559], orgin[1495], orgin[1431], orgin[1367], orgin[1303]} 	= reorder[599:595];
    assign {orgin[280], orgin[216], orgin[152], orgin[88], orgin[24]} 	= reorder[604:600];
    assign {orgin[600], orgin[536], orgin[472], orgin[408], orgin[344]} 	= reorder[609:605];
    assign {orgin[920], orgin[856], orgin[792], orgin[728], orgin[664]} 	= reorder[614:610];
    assign {orgin[1240], orgin[1176], orgin[1112], orgin[1048], orgin[984]} 	= reorder[619:615];
    assign {orgin[1560], orgin[1496], orgin[1432], orgin[1368], orgin[1304]} 	= reorder[624:620];
    assign {orgin[281], orgin[217], orgin[153], orgin[89], orgin[25]} 	= reorder[629:625];
    assign {orgin[601], orgin[537], orgin[473], orgin[409], orgin[345]} 	= reorder[634:630];
    assign {orgin[921], orgin[857], orgin[793], orgin[729], orgin[665]} 	= reorder[639:635];
    assign {orgin[1241], orgin[1177], orgin[1113], orgin[1049], orgin[985]} 	= reorder[644:640];
    assign {orgin[1561], orgin[1497], orgin[1433], orgin[1369], orgin[1305]} 	= reorder[649:645];
    assign {orgin[282], orgin[218], orgin[154], orgin[90], orgin[26]} 	= reorder[654:650];
    assign {orgin[602], orgin[538], orgin[474], orgin[410], orgin[346]} 	= reorder[659:655];
    assign {orgin[922], orgin[858], orgin[794], orgin[730], orgin[666]} 	= reorder[664:660];
    assign {orgin[1242], orgin[1178], orgin[1114], orgin[1050], orgin[986]} 	= reorder[669:665];
    assign {orgin[1562], orgin[1498], orgin[1434], orgin[1370], orgin[1306]} 	= reorder[674:670];
    assign {orgin[283], orgin[219], orgin[155], orgin[91], orgin[27]} 	= reorder[679:675];
    assign {orgin[603], orgin[539], orgin[475], orgin[411], orgin[347]} 	= reorder[684:680];
    assign {orgin[923], orgin[859], orgin[795], orgin[731], orgin[667]} 	= reorder[689:685];
    assign {orgin[1243], orgin[1179], orgin[1115], orgin[1051], orgin[987]} 	= reorder[694:690];
    assign {orgin[1563], orgin[1499], orgin[1435], orgin[1371], orgin[1307]} 	= reorder[699:695];
    assign {orgin[284], orgin[220], orgin[156], orgin[92], orgin[28]} 	= reorder[704:700];
    assign {orgin[604], orgin[540], orgin[476], orgin[412], orgin[348]} 	= reorder[709:705];
    assign {orgin[924], orgin[860], orgin[796], orgin[732], orgin[668]} 	= reorder[714:710];
    assign {orgin[1244], orgin[1180], orgin[1116], orgin[1052], orgin[988]} 	= reorder[719:715];
    assign {orgin[1564], orgin[1500], orgin[1436], orgin[1372], orgin[1308]} 	= reorder[724:720];
    assign {orgin[285], orgin[221], orgin[157], orgin[93], orgin[29]} 	= reorder[729:725];
    assign {orgin[605], orgin[541], orgin[477], orgin[413], orgin[349]} 	= reorder[734:730];
    assign {orgin[925], orgin[861], orgin[797], orgin[733], orgin[669]} 	= reorder[739:735];
    assign {orgin[1245], orgin[1181], orgin[1117], orgin[1053], orgin[989]} 	= reorder[744:740];
    assign {orgin[1565], orgin[1501], orgin[1437], orgin[1373], orgin[1309]} 	= reorder[749:745];
    assign {orgin[286], orgin[222], orgin[158], orgin[94], orgin[30]} 	= reorder[754:750];
    assign {orgin[606], orgin[542], orgin[478], orgin[414], orgin[350]} 	= reorder[759:755];
    assign {orgin[926], orgin[862], orgin[798], orgin[734], orgin[670]} 	= reorder[764:760];
    assign {orgin[1246], orgin[1182], orgin[1118], orgin[1054], orgin[990]} 	= reorder[769:765];
    assign {orgin[1566], orgin[1502], orgin[1438], orgin[1374], orgin[1310]} 	= reorder[774:770];
    assign {orgin[287], orgin[223], orgin[159], orgin[95], orgin[31]} 	= reorder[779:775];
    assign {orgin[607], orgin[543], orgin[479], orgin[415], orgin[351]} 	= reorder[784:780];
    assign {orgin[927], orgin[863], orgin[799], orgin[735], orgin[671]} 	= reorder[789:785];
    assign {orgin[1247], orgin[1183], orgin[1119], orgin[1055], orgin[991]} 	= reorder[794:790];
    assign {orgin[1567], orgin[1503], orgin[1439], orgin[1375], orgin[1311]} 	= reorder[799:795];
    assign {orgin[288], orgin[224], orgin[160], orgin[96], orgin[32]} 	= reorder[804:800];
    assign {orgin[608], orgin[544], orgin[480], orgin[416], orgin[352]} 	= reorder[809:805];
    assign {orgin[928], orgin[864], orgin[800], orgin[736], orgin[672]} 	= reorder[814:810];
    assign {orgin[1248], orgin[1184], orgin[1120], orgin[1056], orgin[992]} 	= reorder[819:815];
    assign {orgin[1568], orgin[1504], orgin[1440], orgin[1376], orgin[1312]} 	= reorder[824:820];
    assign {orgin[289], orgin[225], orgin[161], orgin[97], orgin[33]} 	= reorder[829:825];
    assign {orgin[609], orgin[545], orgin[481], orgin[417], orgin[353]} 	= reorder[834:830];
    assign {orgin[929], orgin[865], orgin[801], orgin[737], orgin[673]} 	= reorder[839:835];
    assign {orgin[1249], orgin[1185], orgin[1121], orgin[1057], orgin[993]} 	= reorder[844:840];
    assign {orgin[1569], orgin[1505], orgin[1441], orgin[1377], orgin[1313]} 	= reorder[849:845];
    assign {orgin[290], orgin[226], orgin[162], orgin[98], orgin[34]} 	= reorder[854:850];
    assign {orgin[610], orgin[546], orgin[482], orgin[418], orgin[354]} 	= reorder[859:855];
    assign {orgin[930], orgin[866], orgin[802], orgin[738], orgin[674]} 	= reorder[864:860];
    assign {orgin[1250], orgin[1186], orgin[1122], orgin[1058], orgin[994]} 	= reorder[869:865];
    assign {orgin[1570], orgin[1506], orgin[1442], orgin[1378], orgin[1314]} 	= reorder[874:870];
    assign {orgin[291], orgin[227], orgin[163], orgin[99], orgin[35]} 	= reorder[879:875];
    assign {orgin[611], orgin[547], orgin[483], orgin[419], orgin[355]} 	= reorder[884:880];
    assign {orgin[931], orgin[867], orgin[803], orgin[739], orgin[675]} 	= reorder[889:885];
    assign {orgin[1251], orgin[1187], orgin[1123], orgin[1059], orgin[995]} 	= reorder[894:890];
    assign {orgin[1571], orgin[1507], orgin[1443], orgin[1379], orgin[1315]} 	= reorder[899:895];
    assign {orgin[292], orgin[228], orgin[164], orgin[100], orgin[36]} 	= reorder[904:900];
    assign {orgin[612], orgin[548], orgin[484], orgin[420], orgin[356]} 	= reorder[909:905];
    assign {orgin[932], orgin[868], orgin[804], orgin[740], orgin[676]} 	= reorder[914:910];
    assign {orgin[1252], orgin[1188], orgin[1124], orgin[1060], orgin[996]} 	= reorder[919:915];
    assign {orgin[1572], orgin[1508], orgin[1444], orgin[1380], orgin[1316]} 	= reorder[924:920];
    assign {orgin[293], orgin[229], orgin[165], orgin[101], orgin[37]} 	= reorder[929:925];
    assign {orgin[613], orgin[549], orgin[485], orgin[421], orgin[357]} 	= reorder[934:930];
    assign {orgin[933], orgin[869], orgin[805], orgin[741], orgin[677]} 	= reorder[939:935];
    assign {orgin[1253], orgin[1189], orgin[1125], orgin[1061], orgin[997]} 	= reorder[944:940];
    assign {orgin[1573], orgin[1509], orgin[1445], orgin[1381], orgin[1317]} 	= reorder[949:945];
    assign {orgin[294], orgin[230], orgin[166], orgin[102], orgin[38]} 	= reorder[954:950];
    assign {orgin[614], orgin[550], orgin[486], orgin[422], orgin[358]} 	= reorder[959:955];
    assign {orgin[934], orgin[870], orgin[806], orgin[742], orgin[678]} 	= reorder[964:960];
    assign {orgin[1254], orgin[1190], orgin[1126], orgin[1062], orgin[998]} 	= reorder[969:965];
    assign {orgin[1574], orgin[1510], orgin[1446], orgin[1382], orgin[1318]} 	= reorder[974:970];
    assign {orgin[295], orgin[231], orgin[167], orgin[103], orgin[39]} 	= reorder[979:975];
    assign {orgin[615], orgin[551], orgin[487], orgin[423], orgin[359]} 	= reorder[984:980];
    assign {orgin[935], orgin[871], orgin[807], orgin[743], orgin[679]} 	= reorder[989:985];
    assign {orgin[1255], orgin[1191], orgin[1127], orgin[1063], orgin[999]} 	= reorder[994:990];
    assign {orgin[1575], orgin[1511], orgin[1447], orgin[1383], orgin[1319]} 	= reorder[999:995];
    assign {orgin[296], orgin[232], orgin[168], orgin[104], orgin[40]} 	= reorder[1004:1000];
    assign {orgin[616], orgin[552], orgin[488], orgin[424], orgin[360]} 	= reorder[1009:1005];
    assign {orgin[936], orgin[872], orgin[808], orgin[744], orgin[680]} 	= reorder[1014:1010];
    assign {orgin[1256], orgin[1192], orgin[1128], orgin[1064], orgin[1000]} 	= reorder[1019:1015];
    assign {orgin[1576], orgin[1512], orgin[1448], orgin[1384], orgin[1320]} 	= reorder[1024:1020];
    assign {orgin[297], orgin[233], orgin[169], orgin[105], orgin[41]} 	= reorder[1029:1025];
    assign {orgin[617], orgin[553], orgin[489], orgin[425], orgin[361]} 	= reorder[1034:1030];
    assign {orgin[937], orgin[873], orgin[809], orgin[745], orgin[681]} 	= reorder[1039:1035];
    assign {orgin[1257], orgin[1193], orgin[1129], orgin[1065], orgin[1001]} 	= reorder[1044:1040];
    assign {orgin[1577], orgin[1513], orgin[1449], orgin[1385], orgin[1321]} 	= reorder[1049:1045];
    assign {orgin[298], orgin[234], orgin[170], orgin[106], orgin[42]} 	= reorder[1054:1050];
    assign {orgin[618], orgin[554], orgin[490], orgin[426], orgin[362]} 	= reorder[1059:1055];
    assign {orgin[938], orgin[874], orgin[810], orgin[746], orgin[682]} 	= reorder[1064:1060];
    assign {orgin[1258], orgin[1194], orgin[1130], orgin[1066], orgin[1002]} 	= reorder[1069:1065];
    assign {orgin[1578], orgin[1514], orgin[1450], orgin[1386], orgin[1322]} 	= reorder[1074:1070];
    assign {orgin[299], orgin[235], orgin[171], orgin[107], orgin[43]} 	= reorder[1079:1075];
    assign {orgin[619], orgin[555], orgin[491], orgin[427], orgin[363]} 	= reorder[1084:1080];
    assign {orgin[939], orgin[875], orgin[811], orgin[747], orgin[683]} 	= reorder[1089:1085];
    assign {orgin[1259], orgin[1195], orgin[1131], orgin[1067], orgin[1003]} 	= reorder[1094:1090];
    assign {orgin[1579], orgin[1515], orgin[1451], orgin[1387], orgin[1323]} 	= reorder[1099:1095];
    assign {orgin[300], orgin[236], orgin[172], orgin[108], orgin[44]} 	= reorder[1104:1100];
    assign {orgin[620], orgin[556], orgin[492], orgin[428], orgin[364]} 	= reorder[1109:1105];
    assign {orgin[940], orgin[876], orgin[812], orgin[748], orgin[684]} 	= reorder[1114:1110];
    assign {orgin[1260], orgin[1196], orgin[1132], orgin[1068], orgin[1004]} 	= reorder[1119:1115];
    assign {orgin[1580], orgin[1516], orgin[1452], orgin[1388], orgin[1324]} 	= reorder[1124:1120];
    assign {orgin[301], orgin[237], orgin[173], orgin[109], orgin[45]} 	= reorder[1129:1125];
    assign {orgin[621], orgin[557], orgin[493], orgin[429], orgin[365]} 	= reorder[1134:1130];
    assign {orgin[941], orgin[877], orgin[813], orgin[749], orgin[685]} 	= reorder[1139:1135];
    assign {orgin[1261], orgin[1197], orgin[1133], orgin[1069], orgin[1005]} 	= reorder[1144:1140];
    assign {orgin[1581], orgin[1517], orgin[1453], orgin[1389], orgin[1325]} 	= reorder[1149:1145];
    assign {orgin[302], orgin[238], orgin[174], orgin[110], orgin[46]} 	= reorder[1154:1150];
    assign {orgin[622], orgin[558], orgin[494], orgin[430], orgin[366]} 	= reorder[1159:1155];
    assign {orgin[942], orgin[878], orgin[814], orgin[750], orgin[686]} 	= reorder[1164:1160];
    assign {orgin[1262], orgin[1198], orgin[1134], orgin[1070], orgin[1006]} 	= reorder[1169:1165];
    assign {orgin[1582], orgin[1518], orgin[1454], orgin[1390], orgin[1326]} 	= reorder[1174:1170];
    assign {orgin[303], orgin[239], orgin[175], orgin[111], orgin[47]} 	= reorder[1179:1175];
    assign {orgin[623], orgin[559], orgin[495], orgin[431], orgin[367]} 	= reorder[1184:1180];
    assign {orgin[943], orgin[879], orgin[815], orgin[751], orgin[687]} 	= reorder[1189:1185];
    assign {orgin[1263], orgin[1199], orgin[1135], orgin[1071], orgin[1007]} 	= reorder[1194:1190];
    assign {orgin[1583], orgin[1519], orgin[1455], orgin[1391], orgin[1327]} 	= reorder[1199:1195];
    assign {orgin[304], orgin[240], orgin[176], orgin[112], orgin[48]} 	= reorder[1204:1200];
    assign {orgin[624], orgin[560], orgin[496], orgin[432], orgin[368]} 	= reorder[1209:1205];
    assign {orgin[944], orgin[880], orgin[816], orgin[752], orgin[688]} 	= reorder[1214:1210];
    assign {orgin[1264], orgin[1200], orgin[1136], orgin[1072], orgin[1008]} 	= reorder[1219:1215];
    assign {orgin[1584], orgin[1520], orgin[1456], orgin[1392], orgin[1328]} 	= reorder[1224:1220];
    assign {orgin[305], orgin[241], orgin[177], orgin[113], orgin[49]} 	= reorder[1229:1225];
    assign {orgin[625], orgin[561], orgin[497], orgin[433], orgin[369]} 	= reorder[1234:1230];
    assign {orgin[945], orgin[881], orgin[817], orgin[753], orgin[689]} 	= reorder[1239:1235];
    assign {orgin[1265], orgin[1201], orgin[1137], orgin[1073], orgin[1009]} 	= reorder[1244:1240];
    assign {orgin[1585], orgin[1521], orgin[1457], orgin[1393], orgin[1329]} 	= reorder[1249:1245];
    assign {orgin[306], orgin[242], orgin[178], orgin[114], orgin[50]} 	= reorder[1254:1250];
    assign {orgin[626], orgin[562], orgin[498], orgin[434], orgin[370]} 	= reorder[1259:1255];
    assign {orgin[946], orgin[882], orgin[818], orgin[754], orgin[690]} 	= reorder[1264:1260];
    assign {orgin[1266], orgin[1202], orgin[1138], orgin[1074], orgin[1010]} 	= reorder[1269:1265];
    assign {orgin[1586], orgin[1522], orgin[1458], orgin[1394], orgin[1330]} 	= reorder[1274:1270];
    assign {orgin[307], orgin[243], orgin[179], orgin[115], orgin[51]} 	= reorder[1279:1275];
    assign {orgin[627], orgin[563], orgin[499], orgin[435], orgin[371]} 	= reorder[1284:1280];
    assign {orgin[947], orgin[883], orgin[819], orgin[755], orgin[691]} 	= reorder[1289:1285];
    assign {orgin[1267], orgin[1203], orgin[1139], orgin[1075], orgin[1011]} 	= reorder[1294:1290];
    assign {orgin[1587], orgin[1523], orgin[1459], orgin[1395], orgin[1331]} 	= reorder[1299:1295];
    assign {orgin[308], orgin[244], orgin[180], orgin[116], orgin[52]} 	= reorder[1304:1300];
    assign {orgin[628], orgin[564], orgin[500], orgin[436], orgin[372]} 	= reorder[1309:1305];
    assign {orgin[948], orgin[884], orgin[820], orgin[756], orgin[692]} 	= reorder[1314:1310];
    assign {orgin[1268], orgin[1204], orgin[1140], orgin[1076], orgin[1012]} 	= reorder[1319:1315];
    assign {orgin[1588], orgin[1524], orgin[1460], orgin[1396], orgin[1332]} 	= reorder[1324:1320];
    assign {orgin[309], orgin[245], orgin[181], orgin[117], orgin[53]} 	= reorder[1329:1325];
    assign {orgin[629], orgin[565], orgin[501], orgin[437], orgin[373]} 	= reorder[1334:1330];
    assign {orgin[949], orgin[885], orgin[821], orgin[757], orgin[693]} 	= reorder[1339:1335];
    assign {orgin[1269], orgin[1205], orgin[1141], orgin[1077], orgin[1013]} 	= reorder[1344:1340];
    assign {orgin[1589], orgin[1525], orgin[1461], orgin[1397], orgin[1333]} 	= reorder[1349:1345];
    assign {orgin[310], orgin[246], orgin[182], orgin[118], orgin[54]} 	= reorder[1354:1350];
    assign {orgin[630], orgin[566], orgin[502], orgin[438], orgin[374]} 	= reorder[1359:1355];
    assign {orgin[950], orgin[886], orgin[822], orgin[758], orgin[694]} 	= reorder[1364:1360];
    assign {orgin[1270], orgin[1206], orgin[1142], orgin[1078], orgin[1014]} 	= reorder[1369:1365];
    assign {orgin[1590], orgin[1526], orgin[1462], orgin[1398], orgin[1334]} 	= reorder[1374:1370];
    assign {orgin[311], orgin[247], orgin[183], orgin[119], orgin[55]} 	= reorder[1379:1375];
    assign {orgin[631], orgin[567], orgin[503], orgin[439], orgin[375]} 	= reorder[1384:1380];
    assign {orgin[951], orgin[887], orgin[823], orgin[759], orgin[695]} 	= reorder[1389:1385];
    assign {orgin[1271], orgin[1207], orgin[1143], orgin[1079], orgin[1015]} 	= reorder[1394:1390];
    assign {orgin[1591], orgin[1527], orgin[1463], orgin[1399], orgin[1335]} 	= reorder[1399:1395];
    assign {orgin[312], orgin[248], orgin[184], orgin[120], orgin[56]} 	= reorder[1404:1400];
    assign {orgin[632], orgin[568], orgin[504], orgin[440], orgin[376]} 	= reorder[1409:1405];
    assign {orgin[952], orgin[888], orgin[824], orgin[760], orgin[696]} 	= reorder[1414:1410];
    assign {orgin[1272], orgin[1208], orgin[1144], orgin[1080], orgin[1016]} 	= reorder[1419:1415];
    assign {orgin[1592], orgin[1528], orgin[1464], orgin[1400], orgin[1336]} 	= reorder[1424:1420];
    assign {orgin[313], orgin[249], orgin[185], orgin[121], orgin[57]} 	= reorder[1429:1425];
    assign {orgin[633], orgin[569], orgin[505], orgin[441], orgin[377]} 	= reorder[1434:1430];
    assign {orgin[953], orgin[889], orgin[825], orgin[761], orgin[697]} 	= reorder[1439:1435];
    assign {orgin[1273], orgin[1209], orgin[1145], orgin[1081], orgin[1017]} 	= reorder[1444:1440];
    assign {orgin[1593], orgin[1529], orgin[1465], orgin[1401], orgin[1337]} 	= reorder[1449:1445];
    assign {orgin[314], orgin[250], orgin[186], orgin[122], orgin[58]} 	= reorder[1454:1450];
    assign {orgin[634], orgin[570], orgin[506], orgin[442], orgin[378]} 	= reorder[1459:1455];
    assign {orgin[954], orgin[890], orgin[826], orgin[762], orgin[698]} 	= reorder[1464:1460];
    assign {orgin[1274], orgin[1210], orgin[1146], orgin[1082], orgin[1018]} 	= reorder[1469:1465];
    assign {orgin[1594], orgin[1530], orgin[1466], orgin[1402], orgin[1338]} 	= reorder[1474:1470];
    assign {orgin[315], orgin[251], orgin[187], orgin[123], orgin[59]} 	= reorder[1479:1475];
    assign {orgin[635], orgin[571], orgin[507], orgin[443], orgin[379]} 	= reorder[1484:1480];
    assign {orgin[955], orgin[891], orgin[827], orgin[763], orgin[699]} 	= reorder[1489:1485];
    assign {orgin[1275], orgin[1211], orgin[1147], orgin[1083], orgin[1019]} 	= reorder[1494:1490];
    assign {orgin[1595], orgin[1531], orgin[1467], orgin[1403], orgin[1339]} 	= reorder[1499:1495];
    assign {orgin[316], orgin[252], orgin[188], orgin[124], orgin[60]} 	= reorder[1504:1500];
    assign {orgin[636], orgin[572], orgin[508], orgin[444], orgin[380]} 	= reorder[1509:1505];
    assign {orgin[956], orgin[892], orgin[828], orgin[764], orgin[700]} 	= reorder[1514:1510];
    assign {orgin[1276], orgin[1212], orgin[1148], orgin[1084], orgin[1020]} 	= reorder[1519:1515];
    assign {orgin[1596], orgin[1532], orgin[1468], orgin[1404], orgin[1340]} 	= reorder[1524:1520];
    assign {orgin[317], orgin[253], orgin[189], orgin[125], orgin[61]} 	= reorder[1529:1525];
    assign {orgin[637], orgin[573], orgin[509], orgin[445], orgin[381]} 	= reorder[1534:1530];
    assign {orgin[957], orgin[893], orgin[829], orgin[765], orgin[701]} 	= reorder[1539:1535];
    assign {orgin[1277], orgin[1213], orgin[1149], orgin[1085], orgin[1021]} 	= reorder[1544:1540];
    assign {orgin[1597], orgin[1533], orgin[1469], orgin[1405], orgin[1341]} 	= reorder[1549:1545];
    assign {orgin[318], orgin[254], orgin[190], orgin[126], orgin[62]} 	= reorder[1554:1550];
    assign {orgin[638], orgin[574], orgin[510], orgin[446], orgin[382]} 	= reorder[1559:1555];
    assign {orgin[958], orgin[894], orgin[830], orgin[766], orgin[702]} 	= reorder[1564:1560];
    assign {orgin[1278], orgin[1214], orgin[1150], orgin[1086], orgin[1022]} 	= reorder[1569:1565];
    assign {orgin[1598], orgin[1534], orgin[1470], orgin[1406], orgin[1342]} 	= reorder[1574:1570];
    assign {orgin[319], orgin[255], orgin[191], orgin[127], orgin[63]} 	= reorder[1579:1575];
    assign {orgin[639], orgin[575], orgin[511], orgin[447], orgin[383]} 	= reorder[1584:1580];
    assign {orgin[959], orgin[895], orgin[831], orgin[767], orgin[703]} 	= reorder[1589:1585];
    assign {orgin[1279], orgin[1215], orgin[1151], orgin[1087], orgin[1023]} 	= reorder[1594:1590];
    assign {orgin[1599], orgin[1535], orgin[1471], orgin[1407], orgin[1343]} 	= reorder[1599:1595];
endmodule
